module top_module(output one);
assign one = 1;
endmodule
